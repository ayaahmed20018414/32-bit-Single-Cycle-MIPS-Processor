module and_gate(input IN1,input IN2,output OUT);

assign OUT= IN1 & IN2;

endmodule
